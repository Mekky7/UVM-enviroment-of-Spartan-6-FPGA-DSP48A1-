package shared_pkg;
typedef enum  {SHIFT,ROTATE} mode_e;
typedef enum  {RIGHT,LEFT}   direction_e;
bit parameter_comb;    
endpackage